BZh91AY&SY�g� F_�Py���߰����P�ԃjɡT� ��a�i�&��  h���A�ɓ&F�L�LD$�hSM�������  =&����a2dɑ��4�# C �BhM4����Ѡ	�4 ���3X
a+���p*�_GK)41���	 V:!,�,���Y����=֐D~	��3HնZN'��خ��xժ"(E�-��͛����T㰱�(��"��L[�;���م�
��wn�<̀��xѨ�Y�jr����.�w�d*��GU�%�w��+\a7�Q{�m䗭���eW���v��whl��~��X����У �+R�{b��^g|�d�¢���d �"�X�S�3�t�4]�����r��]��눔��k��2s�Γ'_�h{~bb(�fn�f�%�\J<$��6Z�S�Q��19}��)I{��Y��©ʒ�^�.�_M��������
,>�z�H~/ng1c���S:pJ���*�R�msK���&���II��a�RŨ�̩]X�~�6Ph)8�Qա�3���!-�#���Q>�u�ܜ����	�Z�Cz�g��Ԕ!�j�sE�ha�R��R@Z���J���vUi�M�� �%�ϔ�6�0r�!�Ɯ�A���*��	�o8��zr@�8ћ�	7�$7�	�VSB�q*��BhZ�Y�d
�*���e�q���#Mt��W��b�w:zJx�q��p6��3��8+n��T%�x�[�x9��$v�C��jt=7:���	�L�5���װ��O"#N	kJaO#�Qp�(�Aa��9�x�5yKl�0,	�~|��Cc&n"�1K��NN��vS4Bs�i+t��T��!�d&�0Ѝ��w$S�	��